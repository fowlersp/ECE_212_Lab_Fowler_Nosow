//--------------------------------------------------------------
// adder.sv - 32-bit adder
// Dvid_Harris@hmc.edu and Sarah_Harris@hmc.edu 23 October 2005
// Updated to SystemVerilog dmh 12 November 2010
// Refactored into separate files & updated using additional SystemVerilog
// features by John Nestor May 2018
//--------------------------------------------------------------

module adder(
    input  logic [31:0] a, b,
    output logic [31:0] y
    );

    assign y = a + b;
endmodule
